 


class constraint_41;
	rand bit[4:0]a;
	constraint c1{a<20;}
	constraint c2{a%4 == 0;}
endclass
constraint_41 c1;
module test();
	initial
		begin
			repeat(5)
				begin
					c1=new;
					assert(c1.randomize());
					$display("a=%d",c1.a);
				end
		end
endmodule
